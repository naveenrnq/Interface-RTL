module add(
  input [3:0] a,b,
  output [4:0] sum// cout included
);

  assign sum = a + b;

endmodule
